library verilog;
use verilog.vl_types.all;
entity wordle_vlg_vec_tst is
end wordle_vlg_vec_tst;
